class env extends uvm_env;

  `uvm_component_utils(env)
  




endclass
