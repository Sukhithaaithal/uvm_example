class agent extends uvm_agent;

  `uvm_component_utils(agent)

  function new(string name="agent", uvm_component parent = null);
    super.new(name,parent);
  endfunction

endclass
